// niosII_system.v

// Generated using ACDS version 16.1 196

`timescale 1 ps / 1 ps
module niosII_system (
		input  wire        clk_clk,              //            clk.clk
		output wire [7:0]  green_leds_export,    //     green_leds.export
		input  wire [2:0]  keys_export,          //           keys.export
		output wire [17:0] red_leds_export,      //       red_leds.export
		input  wire        reset_reset_n,        //          reset.reset_n
		inout  wire        sd_card_b_SD_cmd,     //        sd_card.b_SD_cmd
		inout  wire        sd_card_b_SD_dat,     //               .b_SD_dat
		inout  wire        sd_card_b_SD_dat3,    //               .b_SD_dat3
		output wire        sd_card_o_SD_clock,   //               .o_SD_clock
		output wire [12:0] sdram_wire_addr,      //     sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,        //               .ba
		output wire        sdram_wire_cas_n,     //               .cas_n
		output wire        sdram_wire_cke,       //               .cke
		output wire        sdram_wire_cs_n,      //               .cs_n
		inout  wire [31:0] sdram_wire_dq,        //               .dq
		output wire [3:0]  sdram_wire_dqm,       //               .dqm
		output wire        sdram_wire_ras_n,     //               .ras_n
		output wire        sdram_wire_we_n,      //               .we_n
		output wire [6:0]  seven_seg_0_export,   //    seven_seg_0.export
		output wire [6:0]  seven_seg_1_export,   //    seven_seg_1.export
		output wire [6:0]  seven_seg_2_export,   //    seven_seg_2.export
		output wire [6:0]  seven_seg_3_export,   //    seven_seg_3.export
		output wire [6:0]  seven_seg_4_export,   //    seven_seg_4.export
		output wire [6:0]  seven_seg_5_export,   //    seven_seg_5.export
		output wire [6:0]  seven_seg_6_export,   //    seven_seg_6.export
		output wire [6:0]  seven_seg_7_export,   //    seven_seg_7.export
		input  wire [17:0] switches_export,      //       switches.export
		output wire        vga_controller_CLK,   // vga_controller.CLK
		output wire        vga_controller_HS,    //               .HS
		output wire        vga_controller_VS,    //               .VS
		output wire        vga_controller_BLANK, //               .BLANK
		output wire        vga_controller_SYNC,  //               .SYNC
		output wire [7:0]  vga_controller_R,     //               .R
		output wire [7:0]  vga_controller_G,     //               .G
		output wire [7:0]  vga_controller_B      //               .B
	);

	wire         dual_clk_fifo_avalon_dc_buffer_source_valid;                        // DUAL_clk_FIFO:stream_out_valid -> VGA_Controller:valid
	wire  [29:0] dual_clk_fifo_avalon_dc_buffer_source_data;                         // DUAL_clk_FIFO:stream_out_data -> VGA_Controller:data
	wire         dual_clk_fifo_avalon_dc_buffer_source_ready;                        // VGA_Controller:ready -> DUAL_clk_FIFO:stream_out_ready
	wire         dual_clk_fifo_avalon_dc_buffer_source_startofpacket;                // DUAL_clk_FIFO:stream_out_startofpacket -> VGA_Controller:startofpacket
	wire         dual_clk_fifo_avalon_dc_buffer_source_endofpacket;                  // DUAL_clk_FIFO:stream_out_endofpacket -> VGA_Controller:endofpacket
	wire         dma_pixel_buffer_avalon_pixel_source_valid;                         // DMA_Pixel_Buffer:stream_valid -> RGB_Resampler:stream_in_valid
	wire  [15:0] dma_pixel_buffer_avalon_pixel_source_data;                          // DMA_Pixel_Buffer:stream_data -> RGB_Resampler:stream_in_data
	wire         dma_pixel_buffer_avalon_pixel_source_ready;                         // RGB_Resampler:stream_in_ready -> DMA_Pixel_Buffer:stream_ready
	wire         dma_pixel_buffer_avalon_pixel_source_startofpacket;                 // DMA_Pixel_Buffer:stream_startofpacket -> RGB_Resampler:stream_in_startofpacket
	wire         dma_pixel_buffer_avalon_pixel_source_endofpacket;                   // DMA_Pixel_Buffer:stream_endofpacket -> RGB_Resampler:stream_in_endofpacket
	wire         rgb_resampler_avalon_rgb_source_valid;                              // RGB_Resampler:stream_out_valid -> Scaler:stream_in_valid
	wire  [29:0] rgb_resampler_avalon_rgb_source_data;                               // RGB_Resampler:stream_out_data -> Scaler:stream_in_data
	wire         rgb_resampler_avalon_rgb_source_ready;                              // Scaler:stream_in_ready -> RGB_Resampler:stream_out_ready
	wire         rgb_resampler_avalon_rgb_source_startofpacket;                      // RGB_Resampler:stream_out_startofpacket -> Scaler:stream_in_startofpacket
	wire         rgb_resampler_avalon_rgb_source_endofpacket;                        // RGB_Resampler:stream_out_endofpacket -> Scaler:stream_in_endofpacket
	wire         video_clk_vga_clk_clk;                                              // Video_clk:vga_clk_clk -> [DUAL_clk_FIFO:clk_stream_out, VGA_Controller:clk, rst_controller_001:clk]
	wire         dma_pixel_buffer_avalon_pixel_dma_master_waitrequest;               // mm_interconnect_0:DMA_Pixel_Buffer_avalon_pixel_dma_master_waitrequest -> DMA_Pixel_Buffer:master_waitrequest
	wire  [15:0] dma_pixel_buffer_avalon_pixel_dma_master_readdata;                  // mm_interconnect_0:DMA_Pixel_Buffer_avalon_pixel_dma_master_readdata -> DMA_Pixel_Buffer:master_readdata
	wire  [31:0] dma_pixel_buffer_avalon_pixel_dma_master_address;                   // DMA_Pixel_Buffer:master_address -> mm_interconnect_0:DMA_Pixel_Buffer_avalon_pixel_dma_master_address
	wire         dma_pixel_buffer_avalon_pixel_dma_master_read;                      // DMA_Pixel_Buffer:master_read -> mm_interconnect_0:DMA_Pixel_Buffer_avalon_pixel_dma_master_read
	wire         dma_pixel_buffer_avalon_pixel_dma_master_readdatavalid;             // mm_interconnect_0:DMA_Pixel_Buffer_avalon_pixel_dma_master_readdatavalid -> DMA_Pixel_Buffer:master_readdatavalid
	wire         dma_pixel_buffer_avalon_pixel_dma_master_lock;                      // DMA_Pixel_Buffer:master_arbiterlock -> mm_interconnect_0:DMA_Pixel_Buffer_avalon_pixel_dma_master_lock
	wire  [31:0] nios2_qsys_0_data_master_readdata;                                  // mm_interconnect_0:nios2_qsys_0_data_master_readdata -> nios2_qsys_0:d_readdata
	wire         nios2_qsys_0_data_master_waitrequest;                               // mm_interconnect_0:nios2_qsys_0_data_master_waitrequest -> nios2_qsys_0:d_waitrequest
	wire         nios2_qsys_0_data_master_debugaccess;                               // nios2_qsys_0:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:nios2_qsys_0_data_master_debugaccess
	wire  [27:0] nios2_qsys_0_data_master_address;                                   // nios2_qsys_0:d_address -> mm_interconnect_0:nios2_qsys_0_data_master_address
	wire   [3:0] nios2_qsys_0_data_master_byteenable;                                // nios2_qsys_0:d_byteenable -> mm_interconnect_0:nios2_qsys_0_data_master_byteenable
	wire         nios2_qsys_0_data_master_read;                                      // nios2_qsys_0:d_read -> mm_interconnect_0:nios2_qsys_0_data_master_read
	wire         nios2_qsys_0_data_master_readdatavalid;                             // mm_interconnect_0:nios2_qsys_0_data_master_readdatavalid -> nios2_qsys_0:d_readdatavalid
	wire         nios2_qsys_0_data_master_write;                                     // nios2_qsys_0:d_write -> mm_interconnect_0:nios2_qsys_0_data_master_write
	wire  [31:0] nios2_qsys_0_data_master_writedata;                                 // nios2_qsys_0:d_writedata -> mm_interconnect_0:nios2_qsys_0_data_master_writedata
	wire  [31:0] nios2_qsys_0_instruction_master_readdata;                           // mm_interconnect_0:nios2_qsys_0_instruction_master_readdata -> nios2_qsys_0:i_readdata
	wire         nios2_qsys_0_instruction_master_waitrequest;                        // mm_interconnect_0:nios2_qsys_0_instruction_master_waitrequest -> nios2_qsys_0:i_waitrequest
	wire  [27:0] nios2_qsys_0_instruction_master_address;                            // nios2_qsys_0:i_address -> mm_interconnect_0:nios2_qsys_0_instruction_master_address
	wire         nios2_qsys_0_instruction_master_read;                               // nios2_qsys_0:i_read -> mm_interconnect_0:nios2_qsys_0_instruction_master_read
	wire         nios2_qsys_0_instruction_master_readdatavalid;                      // mm_interconnect_0:nios2_qsys_0_instruction_master_readdatavalid -> nios2_qsys_0:i_readdatavalid
	wire  [31:0] mm_interconnect_0_dma_pixel_buffer_avalon_control_slave_readdata;   // DMA_Pixel_Buffer:slave_readdata -> mm_interconnect_0:DMA_Pixel_Buffer_avalon_control_slave_readdata
	wire   [1:0] mm_interconnect_0_dma_pixel_buffer_avalon_control_slave_address;    // mm_interconnect_0:DMA_Pixel_Buffer_avalon_control_slave_address -> DMA_Pixel_Buffer:slave_address
	wire         mm_interconnect_0_dma_pixel_buffer_avalon_control_slave_read;       // mm_interconnect_0:DMA_Pixel_Buffer_avalon_control_slave_read -> DMA_Pixel_Buffer:slave_read
	wire   [3:0] mm_interconnect_0_dma_pixel_buffer_avalon_control_slave_byteenable; // mm_interconnect_0:DMA_Pixel_Buffer_avalon_control_slave_byteenable -> DMA_Pixel_Buffer:slave_byteenable
	wire         mm_interconnect_0_dma_pixel_buffer_avalon_control_slave_write;      // mm_interconnect_0:DMA_Pixel_Buffer_avalon_control_slave_write -> DMA_Pixel_Buffer:slave_write
	wire  [31:0] mm_interconnect_0_dma_pixel_buffer_avalon_control_slave_writedata;  // mm_interconnect_0:DMA_Pixel_Buffer_avalon_control_slave_writedata -> DMA_Pixel_Buffer:slave_writedata
	wire  [31:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata;          // nios2_qsys_0:jtag_debug_module_readdata -> mm_interconnect_0:nios2_qsys_0_jtag_debug_module_readdata
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest;       // nios2_qsys_0:jtag_debug_module_waitrequest -> mm_interconnect_0:nios2_qsys_0_jtag_debug_module_waitrequest
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess;       // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_debugaccess -> nios2_qsys_0:jtag_debug_module_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address;           // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_address -> nios2_qsys_0:jtag_debug_module_address
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read;              // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_read -> nios2_qsys_0:jtag_debug_module_read
	wire   [3:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable;        // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_byteenable -> nios2_qsys_0:jtag_debug_module_byteenable
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write;             // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_write -> nios2_qsys_0:jtag_debug_module_write
	wire  [31:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata;         // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_writedata -> nios2_qsys_0:jtag_debug_module_writedata
	wire         mm_interconnect_0_sdram_s1_chipselect;                              // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [31:0] mm_interconnect_0_sdram_s1_readdata;                                // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                             // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_s1_address;                                 // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                                    // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [3:0] mm_interconnect_0_sdram_s1_byteenable;                              // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                           // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                                   // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [31:0] mm_interconnect_0_sdram_s1_writedata;                               // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;         // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;           // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest;        // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;            // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;               // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;              // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;          // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire         mm_interconnect_0_sd_card_avalon_sdcard_slave_chipselect;           // mm_interconnect_0:SD_Card_avalon_sdcard_slave_chipselect -> SD_Card:i_avalon_chip_select
	wire  [31:0] mm_interconnect_0_sd_card_avalon_sdcard_slave_readdata;             // SD_Card:o_avalon_readdata -> mm_interconnect_0:SD_Card_avalon_sdcard_slave_readdata
	wire         mm_interconnect_0_sd_card_avalon_sdcard_slave_waitrequest;          // SD_Card:o_avalon_waitrequest -> mm_interconnect_0:SD_Card_avalon_sdcard_slave_waitrequest
	wire   [7:0] mm_interconnect_0_sd_card_avalon_sdcard_slave_address;              // mm_interconnect_0:SD_Card_avalon_sdcard_slave_address -> SD_Card:i_avalon_address
	wire         mm_interconnect_0_sd_card_avalon_sdcard_slave_read;                 // mm_interconnect_0:SD_Card_avalon_sdcard_slave_read -> SD_Card:i_avalon_read
	wire   [3:0] mm_interconnect_0_sd_card_avalon_sdcard_slave_byteenable;           // mm_interconnect_0:SD_Card_avalon_sdcard_slave_byteenable -> SD_Card:i_avalon_byteenable
	wire         mm_interconnect_0_sd_card_avalon_sdcard_slave_write;                // mm_interconnect_0:SD_Card_avalon_sdcard_slave_write -> SD_Card:i_avalon_write
	wire  [31:0] mm_interconnect_0_sd_card_avalon_sdcard_slave_writedata;            // mm_interconnect_0:SD_Card_avalon_sdcard_slave_writedata -> SD_Card:i_avalon_writedata
	wire  [31:0] mm_interconnect_0_sysid_qsys_0_control_slave_readdata;              // sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_0_control_slave_address;               // mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;                   // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;                     // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire   [9:0] mm_interconnect_0_onchip_memory2_0_s1_address;                      // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;                   // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                        // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;                    // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                        // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire  [31:0] mm_interconnect_0_switches_s1_readdata;                             // switches:readdata -> mm_interconnect_0:switches_s1_readdata
	wire   [1:0] mm_interconnect_0_switches_s1_address;                              // mm_interconnect_0:switches_s1_address -> switches:address
	wire         mm_interconnect_0_red_leds_s1_chipselect;                           // mm_interconnect_0:red_leds_s1_chipselect -> red_leds:chipselect
	wire  [31:0] mm_interconnect_0_red_leds_s1_readdata;                             // red_leds:readdata -> mm_interconnect_0:red_leds_s1_readdata
	wire   [1:0] mm_interconnect_0_red_leds_s1_address;                              // mm_interconnect_0:red_leds_s1_address -> red_leds:address
	wire         mm_interconnect_0_red_leds_s1_write;                                // mm_interconnect_0:red_leds_s1_write -> red_leds:write_n
	wire  [31:0] mm_interconnect_0_red_leds_s1_writedata;                            // mm_interconnect_0:red_leds_s1_writedata -> red_leds:writedata
	wire         mm_interconnect_0_green_leds_s1_chipselect;                         // mm_interconnect_0:green_leds_s1_chipselect -> green_leds:chipselect
	wire  [31:0] mm_interconnect_0_green_leds_s1_readdata;                           // green_leds:readdata -> mm_interconnect_0:green_leds_s1_readdata
	wire   [1:0] mm_interconnect_0_green_leds_s1_address;                            // mm_interconnect_0:green_leds_s1_address -> green_leds:address
	wire         mm_interconnect_0_green_leds_s1_write;                              // mm_interconnect_0:green_leds_s1_write -> green_leds:write_n
	wire  [31:0] mm_interconnect_0_green_leds_s1_writedata;                          // mm_interconnect_0:green_leds_s1_writedata -> green_leds:writedata
	wire         mm_interconnect_0_keys_s1_chipselect;                               // mm_interconnect_0:KEYS_s1_chipselect -> KEYS:chipselect
	wire  [31:0] mm_interconnect_0_keys_s1_readdata;                                 // KEYS:readdata -> mm_interconnect_0:KEYS_s1_readdata
	wire   [1:0] mm_interconnect_0_keys_s1_address;                                  // mm_interconnect_0:KEYS_s1_address -> KEYS:address
	wire         mm_interconnect_0_keys_s1_write;                                    // mm_interconnect_0:KEYS_s1_write -> KEYS:write_n
	wire  [31:0] mm_interconnect_0_keys_s1_writedata;                                // mm_interconnect_0:KEYS_s1_writedata -> KEYS:writedata
	wire         mm_interconnect_0_seven_seg_0_s1_chipselect;                        // mm_interconnect_0:seven_seg_0_s1_chipselect -> seven_seg_0:chipselect
	wire  [31:0] mm_interconnect_0_seven_seg_0_s1_readdata;                          // seven_seg_0:readdata -> mm_interconnect_0:seven_seg_0_s1_readdata
	wire   [1:0] mm_interconnect_0_seven_seg_0_s1_address;                           // mm_interconnect_0:seven_seg_0_s1_address -> seven_seg_0:address
	wire         mm_interconnect_0_seven_seg_0_s1_write;                             // mm_interconnect_0:seven_seg_0_s1_write -> seven_seg_0:write_n
	wire  [31:0] mm_interconnect_0_seven_seg_0_s1_writedata;                         // mm_interconnect_0:seven_seg_0_s1_writedata -> seven_seg_0:writedata
	wire         mm_interconnect_0_seven_seg_1_s1_chipselect;                        // mm_interconnect_0:seven_seg_1_s1_chipselect -> seven_seg_1:chipselect
	wire  [31:0] mm_interconnect_0_seven_seg_1_s1_readdata;                          // seven_seg_1:readdata -> mm_interconnect_0:seven_seg_1_s1_readdata
	wire   [1:0] mm_interconnect_0_seven_seg_1_s1_address;                           // mm_interconnect_0:seven_seg_1_s1_address -> seven_seg_1:address
	wire         mm_interconnect_0_seven_seg_1_s1_write;                             // mm_interconnect_0:seven_seg_1_s1_write -> seven_seg_1:write_n
	wire  [31:0] mm_interconnect_0_seven_seg_1_s1_writedata;                         // mm_interconnect_0:seven_seg_1_s1_writedata -> seven_seg_1:writedata
	wire         mm_interconnect_0_seven_seg_2_s1_chipselect;                        // mm_interconnect_0:seven_seg_2_s1_chipselect -> seven_seg_2:chipselect
	wire  [31:0] mm_interconnect_0_seven_seg_2_s1_readdata;                          // seven_seg_2:readdata -> mm_interconnect_0:seven_seg_2_s1_readdata
	wire   [1:0] mm_interconnect_0_seven_seg_2_s1_address;                           // mm_interconnect_0:seven_seg_2_s1_address -> seven_seg_2:address
	wire         mm_interconnect_0_seven_seg_2_s1_write;                             // mm_interconnect_0:seven_seg_2_s1_write -> seven_seg_2:write_n
	wire  [31:0] mm_interconnect_0_seven_seg_2_s1_writedata;                         // mm_interconnect_0:seven_seg_2_s1_writedata -> seven_seg_2:writedata
	wire         mm_interconnect_0_seven_seg_3_s1_chipselect;                        // mm_interconnect_0:seven_seg_3_s1_chipselect -> seven_seg_3:chipselect
	wire  [31:0] mm_interconnect_0_seven_seg_3_s1_readdata;                          // seven_seg_3:readdata -> mm_interconnect_0:seven_seg_3_s1_readdata
	wire   [1:0] mm_interconnect_0_seven_seg_3_s1_address;                           // mm_interconnect_0:seven_seg_3_s1_address -> seven_seg_3:address
	wire         mm_interconnect_0_seven_seg_3_s1_write;                             // mm_interconnect_0:seven_seg_3_s1_write -> seven_seg_3:write_n
	wire  [31:0] mm_interconnect_0_seven_seg_3_s1_writedata;                         // mm_interconnect_0:seven_seg_3_s1_writedata -> seven_seg_3:writedata
	wire         mm_interconnect_0_seven_seg_4_s1_chipselect;                        // mm_interconnect_0:seven_seg_4_s1_chipselect -> seven_seg_4:chipselect
	wire  [31:0] mm_interconnect_0_seven_seg_4_s1_readdata;                          // seven_seg_4:readdata -> mm_interconnect_0:seven_seg_4_s1_readdata
	wire   [1:0] mm_interconnect_0_seven_seg_4_s1_address;                           // mm_interconnect_0:seven_seg_4_s1_address -> seven_seg_4:address
	wire         mm_interconnect_0_seven_seg_4_s1_write;                             // mm_interconnect_0:seven_seg_4_s1_write -> seven_seg_4:write_n
	wire  [31:0] mm_interconnect_0_seven_seg_4_s1_writedata;                         // mm_interconnect_0:seven_seg_4_s1_writedata -> seven_seg_4:writedata
	wire         mm_interconnect_0_seven_seg_5_s1_chipselect;                        // mm_interconnect_0:seven_seg_5_s1_chipselect -> seven_seg_5:chipselect
	wire  [31:0] mm_interconnect_0_seven_seg_5_s1_readdata;                          // seven_seg_5:readdata -> mm_interconnect_0:seven_seg_5_s1_readdata
	wire   [1:0] mm_interconnect_0_seven_seg_5_s1_address;                           // mm_interconnect_0:seven_seg_5_s1_address -> seven_seg_5:address
	wire         mm_interconnect_0_seven_seg_5_s1_write;                             // mm_interconnect_0:seven_seg_5_s1_write -> seven_seg_5:write_n
	wire  [31:0] mm_interconnect_0_seven_seg_5_s1_writedata;                         // mm_interconnect_0:seven_seg_5_s1_writedata -> seven_seg_5:writedata
	wire         mm_interconnect_0_seven_seg_6_s1_chipselect;                        // mm_interconnect_0:seven_seg_6_s1_chipselect -> seven_seg_6:chipselect
	wire  [31:0] mm_interconnect_0_seven_seg_6_s1_readdata;                          // seven_seg_6:readdata -> mm_interconnect_0:seven_seg_6_s1_readdata
	wire   [1:0] mm_interconnect_0_seven_seg_6_s1_address;                           // mm_interconnect_0:seven_seg_6_s1_address -> seven_seg_6:address
	wire         mm_interconnect_0_seven_seg_6_s1_write;                             // mm_interconnect_0:seven_seg_6_s1_write -> seven_seg_6:write_n
	wire  [31:0] mm_interconnect_0_seven_seg_6_s1_writedata;                         // mm_interconnect_0:seven_seg_6_s1_writedata -> seven_seg_6:writedata
	wire         mm_interconnect_0_system_timer_s1_chipselect;                       // mm_interconnect_0:system_timer_s1_chipselect -> system_timer:chipselect
	wire  [15:0] mm_interconnect_0_system_timer_s1_readdata;                         // system_timer:readdata -> mm_interconnect_0:system_timer_s1_readdata
	wire   [2:0] mm_interconnect_0_system_timer_s1_address;                          // mm_interconnect_0:system_timer_s1_address -> system_timer:address
	wire         mm_interconnect_0_system_timer_s1_write;                            // mm_interconnect_0:system_timer_s1_write -> system_timer:write_n
	wire  [15:0] mm_interconnect_0_system_timer_s1_writedata;                        // mm_interconnect_0:system_timer_s1_writedata -> system_timer:writedata
	wire         mm_interconnect_0_high_res_timer_s1_chipselect;                     // mm_interconnect_0:high_res_timer_s1_chipselect -> high_res_timer:chipselect
	wire  [15:0] mm_interconnect_0_high_res_timer_s1_readdata;                       // high_res_timer:readdata -> mm_interconnect_0:high_res_timer_s1_readdata
	wire   [2:0] mm_interconnect_0_high_res_timer_s1_address;                        // mm_interconnect_0:high_res_timer_s1_address -> high_res_timer:address
	wire         mm_interconnect_0_high_res_timer_s1_write;                          // mm_interconnect_0:high_res_timer_s1_write -> high_res_timer:write_n
	wire  [15:0] mm_interconnect_0_high_res_timer_s1_writedata;                      // mm_interconnect_0:high_res_timer_s1_writedata -> high_res_timer:writedata
	wire         mm_interconnect_0_seven_seg_7_s1_chipselect;                        // mm_interconnect_0:seven_seg_7_s1_chipselect -> seven_seg_7:chipselect
	wire  [31:0] mm_interconnect_0_seven_seg_7_s1_readdata;                          // seven_seg_7:readdata -> mm_interconnect_0:seven_seg_7_s1_readdata
	wire   [1:0] mm_interconnect_0_seven_seg_7_s1_address;                           // mm_interconnect_0:seven_seg_7_s1_address -> seven_seg_7:address
	wire         mm_interconnect_0_seven_seg_7_s1_write;                             // mm_interconnect_0:seven_seg_7_s1_write -> seven_seg_7:write_n
	wire  [31:0] mm_interconnect_0_seven_seg_7_s1_writedata;                         // mm_interconnect_0:seven_seg_7_s1_writedata -> seven_seg_7:writedata
	wire         irq_mapper_receiver0_irq;                                           // KEYS:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                           // system_timer:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                           // high_res_timer:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                           // jtag_uart_0:av_irq -> irq_mapper:receiver3_irq
	wire  [31:0] nios2_qsys_0_d_irq_irq;                                             // irq_mapper:sender_irq -> nios2_qsys_0:d_irq
	wire         scaler_avalon_scaler_source_valid;                                  // Scaler:stream_out_valid -> avalon_st_adapter:in_0_valid
	wire  [29:0] scaler_avalon_scaler_source_data;                                   // Scaler:stream_out_data -> avalon_st_adapter:in_0_data
	wire         scaler_avalon_scaler_source_ready;                                  // avalon_st_adapter:in_0_ready -> Scaler:stream_out_ready
	wire   [1:0] scaler_avalon_scaler_source_channel;                                // Scaler:stream_out_channel -> avalon_st_adapter:in_0_channel
	wire         scaler_avalon_scaler_source_startofpacket;                          // Scaler:stream_out_startofpacket -> avalon_st_adapter:in_0_startofpacket
	wire         scaler_avalon_scaler_source_endofpacket;                            // Scaler:stream_out_endofpacket -> avalon_st_adapter:in_0_endofpacket
	wire         avalon_st_adapter_out_0_valid;                                      // avalon_st_adapter:out_0_valid -> DUAL_clk_FIFO:stream_in_valid
	wire  [29:0] avalon_st_adapter_out_0_data;                                       // avalon_st_adapter:out_0_data -> DUAL_clk_FIFO:stream_in_data
	wire         avalon_st_adapter_out_0_ready;                                      // DUAL_clk_FIFO:stream_in_ready -> avalon_st_adapter:out_0_ready
	wire         avalon_st_adapter_out_0_startofpacket;                              // avalon_st_adapter:out_0_startofpacket -> DUAL_clk_FIFO:stream_in_startofpacket
	wire         avalon_st_adapter_out_0_endofpacket;                                // avalon_st_adapter:out_0_endofpacket -> DUAL_clk_FIFO:stream_in_endofpacket
	wire         rst_controller_reset_out_reset;                                     // rst_controller:reset_out -> [DMA_Pixel_Buffer:reset, DUAL_clk_FIFO:reset_stream_in, KEYS:reset_n, RGB_Resampler:reset, SD_Card:i_reset_n, Scaler:reset, Video_clk:ref_reset_reset, avalon_st_adapter:in_rst_0_reset, green_leds:reset_n, high_res_timer:reset_n, irq_mapper:reset, jtag_uart_0:rst_n, mm_interconnect_0:DMA_Pixel_Buffer_reset_reset_bridge_in_reset_reset, nios2_qsys_0:reset_n, onchip_memory2_0:reset, red_leds:reset_n, rst_translator:in_reset, sdram:reset_n, seven_seg_0:reset_n, seven_seg_1:reset_n, seven_seg_2:reset_n, seven_seg_3:reset_n, seven_seg_4:reset_n, seven_seg_5:reset_n, seven_seg_6:reset_n, seven_seg_7:reset_n, switches:reset_n, sysid_qsys_0:reset_n, system_timer:reset_n]
	wire         rst_controller_reset_out_reset_req;                                 // rst_controller:reset_req -> [nios2_qsys_0:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	wire         nios2_qsys_0_jtag_debug_module_reset_reset;                         // nios2_qsys_0:jtag_debug_module_resetrequest -> [rst_controller:reset_in1, rst_controller_001:reset_in1]
	wire         rst_controller_001_reset_out_reset;                                 // rst_controller_001:reset_out -> [DUAL_clk_FIFO:reset_stream_out, VGA_Controller:reset]

	niosII_system_DMA_Pixel_Buffer dma_pixel_buffer (
		.clk                  (clk_clk),                                                            //                     clk.clk
		.reset                (rst_controller_reset_out_reset),                                     //                   reset.reset
		.master_readdatavalid (dma_pixel_buffer_avalon_pixel_dma_master_readdatavalid),             // avalon_pixel_dma_master.readdatavalid
		.master_waitrequest   (dma_pixel_buffer_avalon_pixel_dma_master_waitrequest),               //                        .waitrequest
		.master_address       (dma_pixel_buffer_avalon_pixel_dma_master_address),                   //                        .address
		.master_arbiterlock   (dma_pixel_buffer_avalon_pixel_dma_master_lock),                      //                        .lock
		.master_read          (dma_pixel_buffer_avalon_pixel_dma_master_read),                      //                        .read
		.master_readdata      (dma_pixel_buffer_avalon_pixel_dma_master_readdata),                  //                        .readdata
		.slave_address        (mm_interconnect_0_dma_pixel_buffer_avalon_control_slave_address),    //    avalon_control_slave.address
		.slave_byteenable     (mm_interconnect_0_dma_pixel_buffer_avalon_control_slave_byteenable), //                        .byteenable
		.slave_read           (mm_interconnect_0_dma_pixel_buffer_avalon_control_slave_read),       //                        .read
		.slave_write          (mm_interconnect_0_dma_pixel_buffer_avalon_control_slave_write),      //                        .write
		.slave_writedata      (mm_interconnect_0_dma_pixel_buffer_avalon_control_slave_writedata),  //                        .writedata
		.slave_readdata       (mm_interconnect_0_dma_pixel_buffer_avalon_control_slave_readdata),   //                        .readdata
		.stream_ready         (dma_pixel_buffer_avalon_pixel_source_ready),                         //     avalon_pixel_source.ready
		.stream_startofpacket (dma_pixel_buffer_avalon_pixel_source_startofpacket),                 //                        .startofpacket
		.stream_endofpacket   (dma_pixel_buffer_avalon_pixel_source_endofpacket),                   //                        .endofpacket
		.stream_valid         (dma_pixel_buffer_avalon_pixel_source_valid),                         //                        .valid
		.stream_data          (dma_pixel_buffer_avalon_pixel_source_data)                           //                        .data
	);

	niosII_system_DUAL_clk_FIFO dual_clk_fifo (
		.clk_stream_in            (clk_clk),                                             //         clock_stream_in.clk
		.reset_stream_in          (rst_controller_reset_out_reset),                      //         reset_stream_in.reset
		.clk_stream_out           (video_clk_vga_clk_clk),                               //        clock_stream_out.clk
		.reset_stream_out         (rst_controller_001_reset_out_reset),                  //        reset_stream_out.reset
		.stream_in_ready          (avalon_st_adapter_out_0_ready),                       //   avalon_dc_buffer_sink.ready
		.stream_in_startofpacket  (avalon_st_adapter_out_0_startofpacket),               //                        .startofpacket
		.stream_in_endofpacket    (avalon_st_adapter_out_0_endofpacket),                 //                        .endofpacket
		.stream_in_valid          (avalon_st_adapter_out_0_valid),                       //                        .valid
		.stream_in_data           (avalon_st_adapter_out_0_data),                        //                        .data
		.stream_out_ready         (dual_clk_fifo_avalon_dc_buffer_source_ready),         // avalon_dc_buffer_source.ready
		.stream_out_startofpacket (dual_clk_fifo_avalon_dc_buffer_source_startofpacket), //                        .startofpacket
		.stream_out_endofpacket   (dual_clk_fifo_avalon_dc_buffer_source_endofpacket),   //                        .endofpacket
		.stream_out_valid         (dual_clk_fifo_avalon_dc_buffer_source_valid),         //                        .valid
		.stream_out_data          (dual_clk_fifo_avalon_dc_buffer_source_data)           //                        .data
	);

	niosII_system_KEYS keys (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_keys_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_keys_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_keys_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_keys_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_keys_s1_readdata),   //                    .readdata
		.in_port    (keys_export),                          // external_connection.export
		.irq        (irq_mapper_receiver0_irq)              //                 irq.irq
	);

	niosII_system_RGB_Resampler rgb_resampler (
		.clk                      (clk_clk),                                            //               clk.clk
		.reset                    (rst_controller_reset_out_reset),                     //             reset.reset
		.stream_in_startofpacket  (dma_pixel_buffer_avalon_pixel_source_startofpacket), //   avalon_rgb_sink.startofpacket
		.stream_in_endofpacket    (dma_pixel_buffer_avalon_pixel_source_endofpacket),   //                  .endofpacket
		.stream_in_valid          (dma_pixel_buffer_avalon_pixel_source_valid),         //                  .valid
		.stream_in_ready          (dma_pixel_buffer_avalon_pixel_source_ready),         //                  .ready
		.stream_in_data           (dma_pixel_buffer_avalon_pixel_source_data),          //                  .data
		.stream_out_ready         (rgb_resampler_avalon_rgb_source_ready),              // avalon_rgb_source.ready
		.stream_out_startofpacket (rgb_resampler_avalon_rgb_source_startofpacket),      //                  .startofpacket
		.stream_out_endofpacket   (rgb_resampler_avalon_rgb_source_endofpacket),        //                  .endofpacket
		.stream_out_valid         (rgb_resampler_avalon_rgb_source_valid),              //                  .valid
		.stream_out_data          (rgb_resampler_avalon_rgb_source_data)                //                  .data
	);

	Altera_UP_SD_Card_Avalon_Interface sd_card (
		.i_avalon_chip_select (mm_interconnect_0_sd_card_avalon_sdcard_slave_chipselect),  // avalon_sdcard_slave.chipselect
		.i_avalon_address     (mm_interconnect_0_sd_card_avalon_sdcard_slave_address),     //                    .address
		.i_avalon_read        (mm_interconnect_0_sd_card_avalon_sdcard_slave_read),        //                    .read
		.i_avalon_write       (mm_interconnect_0_sd_card_avalon_sdcard_slave_write),       //                    .write
		.i_avalon_byteenable  (mm_interconnect_0_sd_card_avalon_sdcard_slave_byteenable),  //                    .byteenable
		.i_avalon_writedata   (mm_interconnect_0_sd_card_avalon_sdcard_slave_writedata),   //                    .writedata
		.o_avalon_readdata    (mm_interconnect_0_sd_card_avalon_sdcard_slave_readdata),    //                    .readdata
		.o_avalon_waitrequest (mm_interconnect_0_sd_card_avalon_sdcard_slave_waitrequest), //                    .waitrequest
		.i_clock              (clk_clk),                                                   //                 clk.clk
		.i_reset_n            (~rst_controller_reset_out_reset),                           //               reset.reset_n
		.b_SD_cmd             (sd_card_b_SD_cmd),                                          //         conduit_end.export
		.b_SD_dat             (sd_card_b_SD_dat),                                          //                    .export
		.b_SD_dat3            (sd_card_b_SD_dat3),                                         //                    .export
		.o_SD_clock           (sd_card_o_SD_clock)                                         //                    .export
	);

	niosII_system_Scaler scaler (
		.clk                      (clk_clk),                                       //                  clk.clk
		.reset                    (rst_controller_reset_out_reset),                //                reset.reset
		.stream_in_startofpacket  (rgb_resampler_avalon_rgb_source_startofpacket), //   avalon_scaler_sink.startofpacket
		.stream_in_endofpacket    (rgb_resampler_avalon_rgb_source_endofpacket),   //                     .endofpacket
		.stream_in_valid          (rgb_resampler_avalon_rgb_source_valid),         //                     .valid
		.stream_in_ready          (rgb_resampler_avalon_rgb_source_ready),         //                     .ready
		.stream_in_data           (rgb_resampler_avalon_rgb_source_data),          //                     .data
		.stream_out_ready         (scaler_avalon_scaler_source_ready),             // avalon_scaler_source.ready
		.stream_out_startofpacket (scaler_avalon_scaler_source_startofpacket),     //                     .startofpacket
		.stream_out_endofpacket   (scaler_avalon_scaler_source_endofpacket),       //                     .endofpacket
		.stream_out_valid         (scaler_avalon_scaler_source_valid),             //                     .valid
		.stream_out_data          (scaler_avalon_scaler_source_data),              //                     .data
		.stream_out_channel       (scaler_avalon_scaler_source_channel)            //                     .channel
	);

	niosII_system_VGA_Controller vga_controller (
		.clk           (video_clk_vga_clk_clk),                               //                clk.clk
		.reset         (rst_controller_001_reset_out_reset),                  //              reset.reset
		.data          (dual_clk_fifo_avalon_dc_buffer_source_data),          //    avalon_vga_sink.data
		.startofpacket (dual_clk_fifo_avalon_dc_buffer_source_startofpacket), //                   .startofpacket
		.endofpacket   (dual_clk_fifo_avalon_dc_buffer_source_endofpacket),   //                   .endofpacket
		.valid         (dual_clk_fifo_avalon_dc_buffer_source_valid),         //                   .valid
		.ready         (dual_clk_fifo_avalon_dc_buffer_source_ready),         //                   .ready
		.VGA_CLK       (vga_controller_CLK),                                  // external_interface.export
		.VGA_HS        (vga_controller_HS),                                   //                   .export
		.VGA_VS        (vga_controller_VS),                                   //                   .export
		.VGA_BLANK     (vga_controller_BLANK),                                //                   .export
		.VGA_SYNC      (vga_controller_SYNC),                                 //                   .export
		.VGA_R         (vga_controller_R),                                    //                   .export
		.VGA_G         (vga_controller_G),                                    //                   .export
		.VGA_B         (vga_controller_B)                                     //                   .export
	);

	niosII_system_Video_clk video_clk (
		.ref_clk_clk        (clk_clk),                        //      ref_clk.clk
		.ref_reset_reset    (rst_controller_reset_out_reset), //    ref_reset.reset
		.vga_clk_clk        (video_clk_vga_clk_clk),          //      vga_clk.clk
		.reset_source_reset ()                                // reset_source.reset
	);

	niosII_system_green_leds green_leds (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_green_leds_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_green_leds_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_green_leds_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_green_leds_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_green_leds_s1_readdata),   //                    .readdata
		.out_port   (green_leds_export)                           // external_connection.export
	);

	niosII_system_high_res_timer high_res_timer (
		.clk        (clk_clk),                                        //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                // reset.reset_n
		.address    (mm_interconnect_0_high_res_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_high_res_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_high_res_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_high_res_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_high_res_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver2_irq)                        //   irq.irq
	);

	niosII_system_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver3_irq)                                     //               irq.irq
	);

	niosII_system_nios2_qsys_0 nios2_qsys_0 (
		.clk                                   (clk_clk),                                                      //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                              //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                           //                          .reset_req
		.d_address                             (nios2_qsys_0_data_master_address),                             //               data_master.address
		.d_byteenable                          (nios2_qsys_0_data_master_byteenable),                          //                          .byteenable
		.d_read                                (nios2_qsys_0_data_master_read),                                //                          .read
		.d_readdata                            (nios2_qsys_0_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (nios2_qsys_0_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (nios2_qsys_0_data_master_write),                               //                          .write
		.d_writedata                           (nios2_qsys_0_data_master_writedata),                           //                          .writedata
		.d_readdatavalid                       (nios2_qsys_0_data_master_readdatavalid),                       //                          .readdatavalid
		.jtag_debug_module_debugaccess_to_roms (nios2_qsys_0_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (nios2_qsys_0_instruction_master_address),                      //        instruction_master.address
		.i_read                                (nios2_qsys_0_instruction_master_read),                         //                          .read
		.i_readdata                            (nios2_qsys_0_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (nios2_qsys_0_instruction_master_waitrequest),                  //                          .waitrequest
		.i_readdatavalid                       (nios2_qsys_0_instruction_master_readdatavalid),                //                          .readdatavalid
		.d_irq                                 (nios2_qsys_0_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios2_qsys_0_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                              // custom_instruction_master.readra
	);

	niosII_system_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),               //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	niosII_system_red_leds red_leds (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_red_leds_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_red_leds_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_red_leds_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_red_leds_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_red_leds_s1_readdata),   //                    .readdata
		.out_port   (red_leds_export)                           // external_connection.export
	);

	niosII_system_sdram sdram (
		.clk            (clk_clk),                                  //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	niosII_system_seven_seg_0 seven_seg_0 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_seven_seg_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_seven_seg_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_seven_seg_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_seven_seg_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_seven_seg_0_s1_readdata),   //                    .readdata
		.out_port   (seven_seg_0_export)                           // external_connection.export
	);

	niosII_system_seven_seg_0 seven_seg_1 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_seven_seg_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_seven_seg_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_seven_seg_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_seven_seg_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_seven_seg_1_s1_readdata),   //                    .readdata
		.out_port   (seven_seg_1_export)                           // external_connection.export
	);

	niosII_system_seven_seg_0 seven_seg_2 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_seven_seg_2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_seven_seg_2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_seven_seg_2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_seven_seg_2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_seven_seg_2_s1_readdata),   //                    .readdata
		.out_port   (seven_seg_2_export)                           // external_connection.export
	);

	niosII_system_seven_seg_0 seven_seg_3 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_seven_seg_3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_seven_seg_3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_seven_seg_3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_seven_seg_3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_seven_seg_3_s1_readdata),   //                    .readdata
		.out_port   (seven_seg_3_export)                           // external_connection.export
	);

	niosII_system_seven_seg_0 seven_seg_4 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_seven_seg_4_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_seven_seg_4_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_seven_seg_4_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_seven_seg_4_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_seven_seg_4_s1_readdata),   //                    .readdata
		.out_port   (seven_seg_4_export)                           // external_connection.export
	);

	niosII_system_seven_seg_0 seven_seg_5 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_seven_seg_5_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_seven_seg_5_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_seven_seg_5_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_seven_seg_5_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_seven_seg_5_s1_readdata),   //                    .readdata
		.out_port   (seven_seg_5_export)                           // external_connection.export
	);

	niosII_system_seven_seg_0 seven_seg_6 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_seven_seg_6_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_seven_seg_6_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_seven_seg_6_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_seven_seg_6_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_seven_seg_6_s1_readdata),   //                    .readdata
		.out_port   (seven_seg_6_export)                           // external_connection.export
	);

	niosII_system_seven_seg_0 seven_seg_7 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_seven_seg_7_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_seven_seg_7_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_seven_seg_7_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_seven_seg_7_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_seven_seg_7_s1_readdata),   //                    .readdata
		.out_port   (seven_seg_7_export)                           // external_connection.export
	);

	niosII_system_switches switches (
		.clk      (clk_clk),                                //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address  (mm_interconnect_0_switches_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_switches_s1_readdata), //                    .readdata
		.in_port  (switches_export)                         // external_connection.export
	);

	niosII_system_sysid_qsys_0 sysid_qsys_0 (
		.clock    (clk_clk),                                               //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                       //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_0_control_slave_address)   //              .address
	);

	niosII_system_system_timer system_timer (
		.clk        (clk_clk),                                      //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              // reset.reset_n
		.address    (mm_interconnect_0_system_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_system_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_system_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_system_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_system_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)                      //   irq.irq
	);

	niosII_system_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                          (clk_clk),                                                            //                                    clk_0_clk.clk
		.DMA_Pixel_Buffer_reset_reset_bridge_in_reset_reset     (rst_controller_reset_out_reset),                                     // DMA_Pixel_Buffer_reset_reset_bridge_in_reset.reset
		.DMA_Pixel_Buffer_avalon_pixel_dma_master_address       (dma_pixel_buffer_avalon_pixel_dma_master_address),                   //     DMA_Pixel_Buffer_avalon_pixel_dma_master.address
		.DMA_Pixel_Buffer_avalon_pixel_dma_master_waitrequest   (dma_pixel_buffer_avalon_pixel_dma_master_waitrequest),               //                                             .waitrequest
		.DMA_Pixel_Buffer_avalon_pixel_dma_master_read          (dma_pixel_buffer_avalon_pixel_dma_master_read),                      //                                             .read
		.DMA_Pixel_Buffer_avalon_pixel_dma_master_readdata      (dma_pixel_buffer_avalon_pixel_dma_master_readdata),                  //                                             .readdata
		.DMA_Pixel_Buffer_avalon_pixel_dma_master_readdatavalid (dma_pixel_buffer_avalon_pixel_dma_master_readdatavalid),             //                                             .readdatavalid
		.DMA_Pixel_Buffer_avalon_pixel_dma_master_lock          (dma_pixel_buffer_avalon_pixel_dma_master_lock),                      //                                             .lock
		.nios2_qsys_0_data_master_address                       (nios2_qsys_0_data_master_address),                                   //                     nios2_qsys_0_data_master.address
		.nios2_qsys_0_data_master_waitrequest                   (nios2_qsys_0_data_master_waitrequest),                               //                                             .waitrequest
		.nios2_qsys_0_data_master_byteenable                    (nios2_qsys_0_data_master_byteenable),                                //                                             .byteenable
		.nios2_qsys_0_data_master_read                          (nios2_qsys_0_data_master_read),                                      //                                             .read
		.nios2_qsys_0_data_master_readdata                      (nios2_qsys_0_data_master_readdata),                                  //                                             .readdata
		.nios2_qsys_0_data_master_readdatavalid                 (nios2_qsys_0_data_master_readdatavalid),                             //                                             .readdatavalid
		.nios2_qsys_0_data_master_write                         (nios2_qsys_0_data_master_write),                                     //                                             .write
		.nios2_qsys_0_data_master_writedata                     (nios2_qsys_0_data_master_writedata),                                 //                                             .writedata
		.nios2_qsys_0_data_master_debugaccess                   (nios2_qsys_0_data_master_debugaccess),                               //                                             .debugaccess
		.nios2_qsys_0_instruction_master_address                (nios2_qsys_0_instruction_master_address),                            //              nios2_qsys_0_instruction_master.address
		.nios2_qsys_0_instruction_master_waitrequest            (nios2_qsys_0_instruction_master_waitrequest),                        //                                             .waitrequest
		.nios2_qsys_0_instruction_master_read                   (nios2_qsys_0_instruction_master_read),                               //                                             .read
		.nios2_qsys_0_instruction_master_readdata               (nios2_qsys_0_instruction_master_readdata),                           //                                             .readdata
		.nios2_qsys_0_instruction_master_readdatavalid          (nios2_qsys_0_instruction_master_readdatavalid),                      //                                             .readdatavalid
		.DMA_Pixel_Buffer_avalon_control_slave_address          (mm_interconnect_0_dma_pixel_buffer_avalon_control_slave_address),    //        DMA_Pixel_Buffer_avalon_control_slave.address
		.DMA_Pixel_Buffer_avalon_control_slave_write            (mm_interconnect_0_dma_pixel_buffer_avalon_control_slave_write),      //                                             .write
		.DMA_Pixel_Buffer_avalon_control_slave_read             (mm_interconnect_0_dma_pixel_buffer_avalon_control_slave_read),       //                                             .read
		.DMA_Pixel_Buffer_avalon_control_slave_readdata         (mm_interconnect_0_dma_pixel_buffer_avalon_control_slave_readdata),   //                                             .readdata
		.DMA_Pixel_Buffer_avalon_control_slave_writedata        (mm_interconnect_0_dma_pixel_buffer_avalon_control_slave_writedata),  //                                             .writedata
		.DMA_Pixel_Buffer_avalon_control_slave_byteenable       (mm_interconnect_0_dma_pixel_buffer_avalon_control_slave_byteenable), //                                             .byteenable
		.green_leds_s1_address                                  (mm_interconnect_0_green_leds_s1_address),                            //                                green_leds_s1.address
		.green_leds_s1_write                                    (mm_interconnect_0_green_leds_s1_write),                              //                                             .write
		.green_leds_s1_readdata                                 (mm_interconnect_0_green_leds_s1_readdata),                           //                                             .readdata
		.green_leds_s1_writedata                                (mm_interconnect_0_green_leds_s1_writedata),                          //                                             .writedata
		.green_leds_s1_chipselect                               (mm_interconnect_0_green_leds_s1_chipselect),                         //                                             .chipselect
		.high_res_timer_s1_address                              (mm_interconnect_0_high_res_timer_s1_address),                        //                            high_res_timer_s1.address
		.high_res_timer_s1_write                                (mm_interconnect_0_high_res_timer_s1_write),                          //                                             .write
		.high_res_timer_s1_readdata                             (mm_interconnect_0_high_res_timer_s1_readdata),                       //                                             .readdata
		.high_res_timer_s1_writedata                            (mm_interconnect_0_high_res_timer_s1_writedata),                      //                                             .writedata
		.high_res_timer_s1_chipselect                           (mm_interconnect_0_high_res_timer_s1_chipselect),                     //                                             .chipselect
		.jtag_uart_0_avalon_jtag_slave_address                  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),            //                jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write                    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),              //                                             .write
		.jtag_uart_0_avalon_jtag_slave_read                     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),               //                                             .read
		.jtag_uart_0_avalon_jtag_slave_readdata                 (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),           //                                             .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata                (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),          //                                             .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest              (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest),        //                                             .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect               (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),         //                                             .chipselect
		.KEYS_s1_address                                        (mm_interconnect_0_keys_s1_address),                                  //                                      KEYS_s1.address
		.KEYS_s1_write                                          (mm_interconnect_0_keys_s1_write),                                    //                                             .write
		.KEYS_s1_readdata                                       (mm_interconnect_0_keys_s1_readdata),                                 //                                             .readdata
		.KEYS_s1_writedata                                      (mm_interconnect_0_keys_s1_writedata),                                //                                             .writedata
		.KEYS_s1_chipselect                                     (mm_interconnect_0_keys_s1_chipselect),                               //                                             .chipselect
		.nios2_qsys_0_jtag_debug_module_address                 (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address),           //               nios2_qsys_0_jtag_debug_module.address
		.nios2_qsys_0_jtag_debug_module_write                   (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write),             //                                             .write
		.nios2_qsys_0_jtag_debug_module_read                    (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read),              //                                             .read
		.nios2_qsys_0_jtag_debug_module_readdata                (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata),          //                                             .readdata
		.nios2_qsys_0_jtag_debug_module_writedata               (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata),         //                                             .writedata
		.nios2_qsys_0_jtag_debug_module_byteenable              (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable),        //                                             .byteenable
		.nios2_qsys_0_jtag_debug_module_waitrequest             (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest),       //                                             .waitrequest
		.nios2_qsys_0_jtag_debug_module_debugaccess             (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess),       //                                             .debugaccess
		.onchip_memory2_0_s1_address                            (mm_interconnect_0_onchip_memory2_0_s1_address),                      //                          onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                              (mm_interconnect_0_onchip_memory2_0_s1_write),                        //                                             .write
		.onchip_memory2_0_s1_readdata                           (mm_interconnect_0_onchip_memory2_0_s1_readdata),                     //                                             .readdata
		.onchip_memory2_0_s1_writedata                          (mm_interconnect_0_onchip_memory2_0_s1_writedata),                    //                                             .writedata
		.onchip_memory2_0_s1_byteenable                         (mm_interconnect_0_onchip_memory2_0_s1_byteenable),                   //                                             .byteenable
		.onchip_memory2_0_s1_chipselect                         (mm_interconnect_0_onchip_memory2_0_s1_chipselect),                   //                                             .chipselect
		.onchip_memory2_0_s1_clken                              (mm_interconnect_0_onchip_memory2_0_s1_clken),                        //                                             .clken
		.red_leds_s1_address                                    (mm_interconnect_0_red_leds_s1_address),                              //                                  red_leds_s1.address
		.red_leds_s1_write                                      (mm_interconnect_0_red_leds_s1_write),                                //                                             .write
		.red_leds_s1_readdata                                   (mm_interconnect_0_red_leds_s1_readdata),                             //                                             .readdata
		.red_leds_s1_writedata                                  (mm_interconnect_0_red_leds_s1_writedata),                            //                                             .writedata
		.red_leds_s1_chipselect                                 (mm_interconnect_0_red_leds_s1_chipselect),                           //                                             .chipselect
		.SD_Card_avalon_sdcard_slave_address                    (mm_interconnect_0_sd_card_avalon_sdcard_slave_address),              //                  SD_Card_avalon_sdcard_slave.address
		.SD_Card_avalon_sdcard_slave_write                      (mm_interconnect_0_sd_card_avalon_sdcard_slave_write),                //                                             .write
		.SD_Card_avalon_sdcard_slave_read                       (mm_interconnect_0_sd_card_avalon_sdcard_slave_read),                 //                                             .read
		.SD_Card_avalon_sdcard_slave_readdata                   (mm_interconnect_0_sd_card_avalon_sdcard_slave_readdata),             //                                             .readdata
		.SD_Card_avalon_sdcard_slave_writedata                  (mm_interconnect_0_sd_card_avalon_sdcard_slave_writedata),            //                                             .writedata
		.SD_Card_avalon_sdcard_slave_byteenable                 (mm_interconnect_0_sd_card_avalon_sdcard_slave_byteenable),           //                                             .byteenable
		.SD_Card_avalon_sdcard_slave_waitrequest                (mm_interconnect_0_sd_card_avalon_sdcard_slave_waitrequest),          //                                             .waitrequest
		.SD_Card_avalon_sdcard_slave_chipselect                 (mm_interconnect_0_sd_card_avalon_sdcard_slave_chipselect),           //                                             .chipselect
		.sdram_s1_address                                       (mm_interconnect_0_sdram_s1_address),                                 //                                     sdram_s1.address
		.sdram_s1_write                                         (mm_interconnect_0_sdram_s1_write),                                   //                                             .write
		.sdram_s1_read                                          (mm_interconnect_0_sdram_s1_read),                                    //                                             .read
		.sdram_s1_readdata                                      (mm_interconnect_0_sdram_s1_readdata),                                //                                             .readdata
		.sdram_s1_writedata                                     (mm_interconnect_0_sdram_s1_writedata),                               //                                             .writedata
		.sdram_s1_byteenable                                    (mm_interconnect_0_sdram_s1_byteenable),                              //                                             .byteenable
		.sdram_s1_readdatavalid                                 (mm_interconnect_0_sdram_s1_readdatavalid),                           //                                             .readdatavalid
		.sdram_s1_waitrequest                                   (mm_interconnect_0_sdram_s1_waitrequest),                             //                                             .waitrequest
		.sdram_s1_chipselect                                    (mm_interconnect_0_sdram_s1_chipselect),                              //                                             .chipselect
		.seven_seg_0_s1_address                                 (mm_interconnect_0_seven_seg_0_s1_address),                           //                               seven_seg_0_s1.address
		.seven_seg_0_s1_write                                   (mm_interconnect_0_seven_seg_0_s1_write),                             //                                             .write
		.seven_seg_0_s1_readdata                                (mm_interconnect_0_seven_seg_0_s1_readdata),                          //                                             .readdata
		.seven_seg_0_s1_writedata                               (mm_interconnect_0_seven_seg_0_s1_writedata),                         //                                             .writedata
		.seven_seg_0_s1_chipselect                              (mm_interconnect_0_seven_seg_0_s1_chipselect),                        //                                             .chipselect
		.seven_seg_1_s1_address                                 (mm_interconnect_0_seven_seg_1_s1_address),                           //                               seven_seg_1_s1.address
		.seven_seg_1_s1_write                                   (mm_interconnect_0_seven_seg_1_s1_write),                             //                                             .write
		.seven_seg_1_s1_readdata                                (mm_interconnect_0_seven_seg_1_s1_readdata),                          //                                             .readdata
		.seven_seg_1_s1_writedata                               (mm_interconnect_0_seven_seg_1_s1_writedata),                         //                                             .writedata
		.seven_seg_1_s1_chipselect                              (mm_interconnect_0_seven_seg_1_s1_chipselect),                        //                                             .chipselect
		.seven_seg_2_s1_address                                 (mm_interconnect_0_seven_seg_2_s1_address),                           //                               seven_seg_2_s1.address
		.seven_seg_2_s1_write                                   (mm_interconnect_0_seven_seg_2_s1_write),                             //                                             .write
		.seven_seg_2_s1_readdata                                (mm_interconnect_0_seven_seg_2_s1_readdata),                          //                                             .readdata
		.seven_seg_2_s1_writedata                               (mm_interconnect_0_seven_seg_2_s1_writedata),                         //                                             .writedata
		.seven_seg_2_s1_chipselect                              (mm_interconnect_0_seven_seg_2_s1_chipselect),                        //                                             .chipselect
		.seven_seg_3_s1_address                                 (mm_interconnect_0_seven_seg_3_s1_address),                           //                               seven_seg_3_s1.address
		.seven_seg_3_s1_write                                   (mm_interconnect_0_seven_seg_3_s1_write),                             //                                             .write
		.seven_seg_3_s1_readdata                                (mm_interconnect_0_seven_seg_3_s1_readdata),                          //                                             .readdata
		.seven_seg_3_s1_writedata                               (mm_interconnect_0_seven_seg_3_s1_writedata),                         //                                             .writedata
		.seven_seg_3_s1_chipselect                              (mm_interconnect_0_seven_seg_3_s1_chipselect),                        //                                             .chipselect
		.seven_seg_4_s1_address                                 (mm_interconnect_0_seven_seg_4_s1_address),                           //                               seven_seg_4_s1.address
		.seven_seg_4_s1_write                                   (mm_interconnect_0_seven_seg_4_s1_write),                             //                                             .write
		.seven_seg_4_s1_readdata                                (mm_interconnect_0_seven_seg_4_s1_readdata),                          //                                             .readdata
		.seven_seg_4_s1_writedata                               (mm_interconnect_0_seven_seg_4_s1_writedata),                         //                                             .writedata
		.seven_seg_4_s1_chipselect                              (mm_interconnect_0_seven_seg_4_s1_chipselect),                        //                                             .chipselect
		.seven_seg_5_s1_address                                 (mm_interconnect_0_seven_seg_5_s1_address),                           //                               seven_seg_5_s1.address
		.seven_seg_5_s1_write                                   (mm_interconnect_0_seven_seg_5_s1_write),                             //                                             .write
		.seven_seg_5_s1_readdata                                (mm_interconnect_0_seven_seg_5_s1_readdata),                          //                                             .readdata
		.seven_seg_5_s1_writedata                               (mm_interconnect_0_seven_seg_5_s1_writedata),                         //                                             .writedata
		.seven_seg_5_s1_chipselect                              (mm_interconnect_0_seven_seg_5_s1_chipselect),                        //                                             .chipselect
		.seven_seg_6_s1_address                                 (mm_interconnect_0_seven_seg_6_s1_address),                           //                               seven_seg_6_s1.address
		.seven_seg_6_s1_write                                   (mm_interconnect_0_seven_seg_6_s1_write),                             //                                             .write
		.seven_seg_6_s1_readdata                                (mm_interconnect_0_seven_seg_6_s1_readdata),                          //                                             .readdata
		.seven_seg_6_s1_writedata                               (mm_interconnect_0_seven_seg_6_s1_writedata),                         //                                             .writedata
		.seven_seg_6_s1_chipselect                              (mm_interconnect_0_seven_seg_6_s1_chipselect),                        //                                             .chipselect
		.seven_seg_7_s1_address                                 (mm_interconnect_0_seven_seg_7_s1_address),                           //                               seven_seg_7_s1.address
		.seven_seg_7_s1_write                                   (mm_interconnect_0_seven_seg_7_s1_write),                             //                                             .write
		.seven_seg_7_s1_readdata                                (mm_interconnect_0_seven_seg_7_s1_readdata),                          //                                             .readdata
		.seven_seg_7_s1_writedata                               (mm_interconnect_0_seven_seg_7_s1_writedata),                         //                                             .writedata
		.seven_seg_7_s1_chipselect                              (mm_interconnect_0_seven_seg_7_s1_chipselect),                        //                                             .chipselect
		.switches_s1_address                                    (mm_interconnect_0_switches_s1_address),                              //                                  switches_s1.address
		.switches_s1_readdata                                   (mm_interconnect_0_switches_s1_readdata),                             //                                             .readdata
		.sysid_qsys_0_control_slave_address                     (mm_interconnect_0_sysid_qsys_0_control_slave_address),               //                   sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata                    (mm_interconnect_0_sysid_qsys_0_control_slave_readdata),              //                                             .readdata
		.system_timer_s1_address                                (mm_interconnect_0_system_timer_s1_address),                          //                              system_timer_s1.address
		.system_timer_s1_write                                  (mm_interconnect_0_system_timer_s1_write),                            //                                             .write
		.system_timer_s1_readdata                               (mm_interconnect_0_system_timer_s1_readdata),                         //                                             .readdata
		.system_timer_s1_writedata                              (mm_interconnect_0_system_timer_s1_writedata),                        //                                             .writedata
		.system_timer_s1_chipselect                             (mm_interconnect_0_system_timer_s1_chipselect)                        //                                             .chipselect
	);

	niosII_system_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.sender_irq    (nios2_qsys_0_d_irq_irq)          //    sender.irq
	);

	niosII_system_avalon_st_adapter #(
		.inBitsPerSymbol (10),
		.inUsePackets    (1),
		.inDataWidth     (30),
		.inChannelWidth  (2),
		.inErrorWidth    (0),
		.inUseEmptyPort  (0),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (0),
		.outDataWidth    (30),
		.outChannelWidth (0),
		.outErrorWidth   (0),
		.outUseEmptyPort (0),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter (
		.in_clk_0_clk        (clk_clk),                                   // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_reset_out_reset),            // in_rst_0.reset
		.in_0_data           (scaler_avalon_scaler_source_data),          //     in_0.data
		.in_0_valid          (scaler_avalon_scaler_source_valid),         //         .valid
		.in_0_ready          (scaler_avalon_scaler_source_ready),         //         .ready
		.in_0_startofpacket  (scaler_avalon_scaler_source_startofpacket), //         .startofpacket
		.in_0_endofpacket    (scaler_avalon_scaler_source_endofpacket),   //         .endofpacket
		.in_0_channel        (scaler_avalon_scaler_source_channel),       //         .channel
		.out_0_data          (avalon_st_adapter_out_0_data),              //    out_0.data
		.out_0_valid         (avalon_st_adapter_out_0_valid),             //         .valid
		.out_0_ready         (avalon_st_adapter_out_0_ready),             //         .ready
		.out_0_startofpacket (avalon_st_adapter_out_0_startofpacket),     //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_out_0_endofpacket)        //         .endofpacket
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                             // reset_in0.reset
		.reset_in1      (nios2_qsys_0_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk            (clk_clk),                                    //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),             // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),         //          .reset_req
		.reset_req_in0  (1'b0),                                       // (terminated)
		.reset_req_in1  (1'b0),                                       // (terminated)
		.reset_in2      (1'b0),                                       // (terminated)
		.reset_req_in2  (1'b0),                                       // (terminated)
		.reset_in3      (1'b0),                                       // (terminated)
		.reset_req_in3  (1'b0),                                       // (terminated)
		.reset_in4      (1'b0),                                       // (terminated)
		.reset_req_in4  (1'b0),                                       // (terminated)
		.reset_in5      (1'b0),                                       // (terminated)
		.reset_req_in5  (1'b0),                                       // (terminated)
		.reset_in6      (1'b0),                                       // (terminated)
		.reset_req_in6  (1'b0),                                       // (terminated)
		.reset_in7      (1'b0),                                       // (terminated)
		.reset_req_in7  (1'b0),                                       // (terminated)
		.reset_in8      (1'b0),                                       // (terminated)
		.reset_req_in8  (1'b0),                                       // (terminated)
		.reset_in9      (1'b0),                                       // (terminated)
		.reset_req_in9  (1'b0),                                       // (terminated)
		.reset_in10     (1'b0),                                       // (terminated)
		.reset_req_in10 (1'b0),                                       // (terminated)
		.reset_in11     (1'b0),                                       // (terminated)
		.reset_req_in11 (1'b0),                                       // (terminated)
		.reset_in12     (1'b0),                                       // (terminated)
		.reset_req_in12 (1'b0),                                       // (terminated)
		.reset_in13     (1'b0),                                       // (terminated)
		.reset_req_in13 (1'b0),                                       // (terminated)
		.reset_in14     (1'b0),                                       // (terminated)
		.reset_req_in14 (1'b0),                                       // (terminated)
		.reset_in15     (1'b0),                                       // (terminated)
		.reset_req_in15 (1'b0)                                        // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                             // reset_in0.reset
		.reset_in1      (nios2_qsys_0_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk            (video_clk_vga_clk_clk),                      //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),         // reset_out.reset
		.reset_req      (),                                           // (terminated)
		.reset_req_in0  (1'b0),                                       // (terminated)
		.reset_req_in1  (1'b0),                                       // (terminated)
		.reset_in2      (1'b0),                                       // (terminated)
		.reset_req_in2  (1'b0),                                       // (terminated)
		.reset_in3      (1'b0),                                       // (terminated)
		.reset_req_in3  (1'b0),                                       // (terminated)
		.reset_in4      (1'b0),                                       // (terminated)
		.reset_req_in4  (1'b0),                                       // (terminated)
		.reset_in5      (1'b0),                                       // (terminated)
		.reset_req_in5  (1'b0),                                       // (terminated)
		.reset_in6      (1'b0),                                       // (terminated)
		.reset_req_in6  (1'b0),                                       // (terminated)
		.reset_in7      (1'b0),                                       // (terminated)
		.reset_req_in7  (1'b0),                                       // (terminated)
		.reset_in8      (1'b0),                                       // (terminated)
		.reset_req_in8  (1'b0),                                       // (terminated)
		.reset_in9      (1'b0),                                       // (terminated)
		.reset_req_in9  (1'b0),                                       // (terminated)
		.reset_in10     (1'b0),                                       // (terminated)
		.reset_req_in10 (1'b0),                                       // (terminated)
		.reset_in11     (1'b0),                                       // (terminated)
		.reset_req_in11 (1'b0),                                       // (terminated)
		.reset_in12     (1'b0),                                       // (terminated)
		.reset_req_in12 (1'b0),                                       // (terminated)
		.reset_in13     (1'b0),                                       // (terminated)
		.reset_req_in13 (1'b0),                                       // (terminated)
		.reset_in14     (1'b0),                                       // (terminated)
		.reset_req_in14 (1'b0),                                       // (terminated)
		.reset_in15     (1'b0),                                       // (terminated)
		.reset_req_in15 (1'b0)                                        // (terminated)
	);

endmodule
